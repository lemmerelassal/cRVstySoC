library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_unsigned.all;

entity fsm is
port (
	
	rst, clk: STD_LOGIC;
	input0, input1, input2, input3, input4, input5, input6, input7: in STD_LOGIC_VECTOR(31 downto 0);
	output0, output1 : out STD_LOGIC_VECTOR(31 downto 0);
mem_rdata : in std_logic_vector(31 downto 0);
mem_wdata, mem_addr : out std_logic_vector(31 downto 0);
mem_re, mem_we : out std_logic;
mem_wack, mem_rdy : in std_logic;
mem_width : out std_logic_vector(1 downto 0)
);
end fsm;

architecture Behavioural of fsm is
signal i_mem_addr, n_mem_addr, i_mem_wdata, n_mem_wdata, pc, n_pc, reg1, n_reg1, reg2, n_reg2, reg6, n_reg6, reg8, n_reg8, reg9, n_reg9, reg10, n_reg10, reg11, n_reg11, reg12, n_reg12, reg13, n_reg13, reg14, n_reg14, reg15, n_reg15, reg16, n_reg16, reg17, n_reg17, reg18, n_reg18, reg19, n_reg19, reg20, n_reg20, reg21, n_reg21, reg22, n_reg22, reg23, n_reg23, reg24, n_reg24, reg25, n_reg25, reg26, n_reg26, reg27, n_reg27, reg28, n_reg28 : STD_LOGIC_VECTOR(31 downto 0);

begin

mem_addr <= i_mem_addr;
mem_wdata <= i_mem_wdata;

process(rst,clk)
begin
	if rst = '1' then
		reg1 <= (others => '0');
		reg2 <= (others => '0');
		reg6 <= (others => '0');
		reg8 <= (others => '0');
		reg9 <= (others => '0');
		reg10 <= (others => '0');
		reg11 <= (others => '0');
		reg12 <= (others => '0');
		reg13 <= (others => '0');
		reg14 <= (others => '0');
		reg15 <= (others => '0');
		reg16 <= (others => '0');
		reg17 <= (others => '0');
		reg18 <= (others => '0');
		reg19 <= (others => '0');
		reg20 <= (others => '0');
		reg21 <= (others => '0');
		reg22 <= (others => '0');
		reg23 <= (others => '0');
		reg24 <= (others => '0');
		reg25 <= (others => '0');
		reg26 <= (others => '0');
		reg27 <= (others => '0');
		reg28 <= (others => '0');
		i_mem_addr <= (others => '0');
		i_mem_wdata <= (others => '0');
		pc <= X"80000000";
	elsif rising_edge(clk) then
		reg1 <= n_reg1;
		reg2 <= n_reg2;
		reg6 <= n_reg6;
		reg8 <= n_reg8;
		reg9 <= n_reg9;
		reg10 <= n_reg10;
		reg11 <= n_reg11;
		reg12 <= n_reg12;
		reg13 <= n_reg13;
		reg14 <= n_reg14;
		reg15 <= n_reg15;
		reg16 <= n_reg16;
		reg17 <= n_reg17;
		reg18 <= n_reg18;
		reg19 <= n_reg19;
		reg20 <= n_reg20;
		reg21 <= n_reg21;
		reg22 <= n_reg22;
		reg23 <= n_reg23;
		reg24 <= n_reg24;
		reg25 <= n_reg25;
		reg26 <= n_reg26;
		reg27 <= n_reg27;
		reg28 <= n_reg28;
		i_mem_addr <= n_mem_addr;
		i_mem_wdata <= n_mem_wdata;
		pc <= n_pc;
	end if;
end process;

process(pc, mem_rdata, mem_rdy, mem_wack, i_mem_addr, i_mem_wdata, reg1, reg2, reg6, reg8, reg9, reg10, reg11, reg12, reg13, reg14, reg15, reg16, reg17, reg18, reg19, reg20, reg21, reg22, reg23, reg24, reg25, reg26, reg27, reg28)
begin
	n_mem_addr <= i_mem_addr;
	n_mem_wdata <= i_mem_wdata;
	mem_re <= '0';
	mem_we <= '0';
	mem_width <= "00";
	n_pc <= pc;
	n_reg1 <= reg1;
	n_reg2 <= reg2;
	n_reg6 <= reg6;
	n_reg8 <= reg8;
	n_reg9 <= reg9;
	n_reg10 <= reg10;
	n_reg11 <= reg11;
	n_reg12 <= reg12;
	n_reg13 <= reg13;
	n_reg14 <= reg14;
	n_reg15 <= reg15;
	n_reg16 <= reg16;
	n_reg17 <= reg17;
	n_reg18 <= reg18;
	n_reg19 <= reg19;
	n_reg20 <= reg20;
	n_reg21 <= reg21;
	n_reg22 <= reg22;
	n_reg23 <= reg23;
	n_reg24 <= reg24;
	n_reg25 <= reg25;
	n_reg26 <= reg26;
	n_reg27 <= reg27;
	n_reg28 <= reg28;
case pc is
	when X"80000800" => n_pc <= X"80000804"; 
 n_reg2 <= X"80000800";

	when X"80000804" => n_pc <= X"80000808"; 
 n_reg2 <= reg2;

	when X"80000808" => 
 n_pc <= X"80000854";

	when X"8000080c" => n_pc <= X"80000810"; 
 n_reg15 <= reg10;

	when X"80000810" => n_pc <= X"80000814"; 
 n_reg10 <= X"00000000";

	when X"80000814" => n_pc <= X"80000818"; 
 if signed(reg11) < signed(reg15) then n_pc <= X"8000081c"; end if;

	when X"80000818" => 
 n_pc <= reg1;

	when X"8000081c" => n_pc <= X"80000820"; 
 n_reg15 <= reg15 - reg11;

	when X"80000820" => n_pc <= X"80000824"; 
 n_reg10 <= reg10 + X"00000001";

	when X"80000824" => 
 n_pc <= X"80000814";

	when X"80000828" => n_pc <= X"8000082c"; 
 if signed(reg11) < signed(reg10) then n_pc <= X"80000830"; end if;

	when X"8000082c" => 
 n_pc <= reg1;

	when X"80000830" => n_pc <= X"80000834"; 
 n_reg10 <= reg10 - reg11;

	when X"80000834" => 
 n_pc <= X"80000828";

	when X"80000838" => n_pc <= X"8000083c"; 
 n_reg14 <= X"00001000";

	when X"8000083c" => n_mem_addr <= reg14; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000840"; n_reg15 <= (others => '0');n_reg15(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000840" => n_pc <= X"80000844"; 
 n_reg15 <= reg15 and X"00000001";

	when X"80000844" => n_pc <= X"80000848"; 
 if signed(reg15) /= X"00000000" then n_pc <= X"8000083c"; end if;

	when X"80000848" => n_pc <= X"8000084c"; 
 n_reg15 <= X"eadbb000";

	when X"8000084c" => mem_width <= "00"; n_mem_addr <= reg15 + X"00000b01"; n_mem_wdata <= reg10; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000850";
 end if;
	when X"80000850" => 
 n_pc <= reg1;

	when X"80000854" => n_pc <= X"80000858"; 
 n_reg10 <= X"80000000";

	when X"80000858" => n_pc <= X"8000085c"; 
 n_reg10 <= reg10;

	when X"8000085c" => 
 n_pc <= X"80001278";

	when X"80000860" => n_pc <= X"80000864"; 
 if unsigned(reg12) >= unsigned(reg13) then n_pc <= X"8000086c"; end if;

	when X"80000864" => n_pc <= X"80000868"; 
 n_reg11 <= reg11 + reg12;

	when X"80000868" => mem_width <= "00"; n_mem_addr <= reg11; n_mem_wdata <= reg10; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000086C";
 end if;
	when X"8000086c" => 
 n_pc <= reg1;

	when X"80000870" => 
 n_pc <= reg1;

	when X"80000874" => n_pc <= X"80000878"; 
 n_reg2 <= reg2 + X"ffffff90";

	when X"80000878" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000068"; n_mem_wdata <= reg8; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000087C";
 end if;
	when X"8000087c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000064"; n_mem_wdata <= reg9; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000880";
 end if;
	when X"80000880" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000060"; n_mem_wdata <= reg18; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000884";
 end if;
	when X"80000884" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000058"; n_mem_wdata <= reg20; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000888";
 end if;
	when X"80000888" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000054"; n_mem_wdata <= reg21; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000088C";
 end if;
	when X"8000088c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000050"; n_mem_wdata <= reg22; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000890";
 end if;
	when X"80000890" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000048"; n_mem_wdata <= reg24; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000894";
 end if;
	when X"80000894" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000040"; n_mem_wdata <= reg26; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000898";
 end if;
	when X"80000898" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000006c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000089C";
 end if;
	when X"8000089c" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000005c"; n_mem_wdata <= reg19; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800008A0";
 end if;
	when X"800008a0" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000004c"; n_mem_wdata <= reg23; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800008A4";
 end if;
	when X"800008a4" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000044"; n_mem_wdata <= reg25; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800008A8";
 end if;
	when X"800008a8" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg27; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800008AC";
 end if;
	when X"800008ac" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000008"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800008B0";
 end if;
	when X"800008b0" => n_pc <= X"800008b4"; 

 n_reg21 <= reg11;

	when X"800008b4" => n_mem_addr <= reg2 + X"00000070"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800008B8"; n_reg26 <= (others => '0');n_reg26(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800008b8" => n_mem_addr <= reg2 + X"00000074"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800008BC"; n_reg9 <= (others => '0');n_reg9(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800008bc" => n_pc <= X"800008c0"; 
 n_reg20 <= reg10;

	when X"800008c0" => n_pc <= X"800008c4"; 
 n_reg18 <= reg12;

	when X"800008c4" => n_pc <= X"800008c8"; 
 n_reg22 <= reg13;

	when X"800008c8" => n_pc <= X"800008cc"; 
 n_reg8 <= reg14;

	when X"800008cc" => n_pc <= X"800008d0"; 
 n_reg11 <= reg16;

	when X"800008d0" => n_pc <= X"800008d4"; 
 n_reg24 <= reg17;

	when X"800008d4" => n_pc <= X"800008d8"; 
 if signed(reg14) /= X"00000000" then n_pc <= X"800008dc"; end if;

	when X"800008d8" => n_pc <= X"800008dc"; 
 n_reg9 <= reg9 and X"ffffffef";

	when X"800008dc" => n_pc <= X"800008e0"; 
 n_reg25 <= reg9 and X"00000400";

	when X"800008e0" => n_pc <= X"800008e4"; 
 if signed(reg25) = X"00000000" then n_pc <= X"800008e8"; end if;

	when X"800008e4" => n_pc <= X"800008e8"; 
 if signed(reg8) = X"00000000" then n_pc <= X"80000954"; end if;

	when X"800008e8" => n_pc <= X"800008ec"; 
 n_reg14 <= reg9 and X"00000020";

	when X"800008ec" => n_pc <= X"800008f0"; 
 n_reg19 <= X"00000061";

	when X"800008f0" => n_pc <= X"800008f4"; 
 if signed(reg14) = X"00000000" then n_pc <= X"800008f8"; end if;

	when X"800008f4" => n_pc <= X"800008f8"; 
 n_reg19 <= X"00000041";

	when X"800008f8" => n_pc <= X"800008fc"; 
 n_reg23 <= reg8;

	when X"800008fc" => n_pc <= X"80000900"; 
 n_reg27 <= reg2 + X"00000010";

	when X"80000900" => n_pc <= X"80000904"; 
 n_reg8 <= X"00000000";

	when X"80000904" => n_pc <= X"80000908"; 
 n_reg19 <= reg19 + X"fffffff6";

	when X"80000908" => n_pc <= X"8000090c"; 
 n_reg10 <= reg23;

	when X"8000090c" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg11; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000910";
 end if;
	when X"80000910" => 
 n_reg1 <= X"80000914"; n_pc <= X"80000828";

	when X"80000914" => n_pc <= X"80000918"; 
 n_reg15 <= X"00000009";

	when X"80000918" => n_mem_addr <= reg2 + X"0000000c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"8000091C"; n_reg11 <= (others => '0');n_reg11(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"8000091c" => n_pc <= X"80000920"; 
 n_reg14 <= reg10 and X"000000ff";

	when X"80000920" => n_pc <= X"80000924"; 
 if unsigned(reg15) < unsigned(reg10) then n_pc <= X"80000990"; end if;

	when X"80000924" => n_pc <= X"80000928"; 
 n_reg14 <= reg14 + X"00000030";

	when X"80000928" => n_pc <= X"8000092c"; 
 n_reg14 <= reg14 and X"000000ff";

	when X"8000092c" => n_pc <= X"80000930"; 
 n_reg10 <= reg23;

	when X"80000930" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg11; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000934";
 end if;
	when X"80000934" => mem_width <= "00"; n_mem_addr <= reg27; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000938";
 end if;
	when X"80000938" => 
 n_reg1 <= X"8000093C"; n_pc <= X"8000080c";

	when X"8000093c" => n_mem_addr <= reg2 + X"0000000c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000940"; n_reg11 <= (others => '0');n_reg11(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000940" => n_pc <= X"80000944"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000944" => n_pc <= X"80000948"; 
 if unsigned(reg23) < unsigned(reg11) then n_pc <= X"80000954"; end if;

	when X"80000948" => n_pc <= X"8000094c"; 
 n_reg15 <= X"00000020";

	when X"8000094c" => n_pc <= X"80000950"; 
 n_reg27 <= reg27 + X"00000001";

	when X"80000950" => n_pc <= X"80000954"; 
 if signed(reg8) /= signed(reg15) then n_pc <= X"80000988"; end if;

	when X"80000954" => n_pc <= X"80000958"; 
 n_reg19 <= reg9 and X"00000002";

	when X"80000958" => n_pc <= X"8000095c"; 
 if signed(reg19) /= X"00000000" then n_pc <= X"800009c4"; end if;

	when X"8000095c" => n_pc <= X"80000960"; 
 n_reg14 <= reg9 and X"00000001";

	when X"80000960" => n_pc <= X"80000964"; 
 if signed(reg26) = X"00000000" then n_pc <= X"8000097c"; end if;

	when X"80000964" => n_pc <= X"80000968"; 
 if signed(reg14) = X"00000000" then n_pc <= X"8000097c"; end if;

	when X"80000968" => n_mem_addr <= reg2 + X"00000008"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"8000096C"; n_reg15 <= (others => '0');n_reg15(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"8000096c" => n_pc <= X"80000970"; 
 if signed(reg15) /= X"00000000" then n_pc <= X"80000978"; end if;

	when X"80000970" => n_pc <= X"80000974"; 
 n_reg13 <= reg9 and X"0000000c";

	when X"80000974" => n_pc <= X"80000978"; 
 if signed(reg13) = X"00000000" then n_pc <= X"8000097c"; end if;

	when X"80000978" => n_pc <= X"8000097c"; 
 n_reg26 <= reg26 + X"ffffffff";


	when X"8000097c" => n_pc <= X"80000980"; 
 n_reg13 <= X"00000020";

	when X"80000980" => n_pc <= X"80000984"; 
 n_reg12 <= X"00000030";

	when X"80000984" => 
 n_pc <= X"800009a8";

	when X"80000988" => n_pc <= X"8000098c"; 
 n_reg23 <= reg10;

	when X"8000098c" => 
 n_pc <= X"80000908";

	when X"80000990" => n_pc <= X"80000994"; 
 n_reg14 <= reg14 + reg19;

	when X"80000994" => 
 n_pc <= X"80000928";

	when X"80000998" => n_pc <= X"8000099c"; 
 n_reg15 <= reg2 + X"00000010";

	when X"8000099c" => n_pc <= X"800009a0"; 
 n_reg10 <= reg15 + reg8;

	when X"800009a0" => mem_width <= "00"; n_mem_addr <= reg10; n_mem_wdata <= reg12; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800009A4";
 end if;
	when X"800009a4" => n_pc <= X"800009a8"; 
 n_reg8 <= reg8 + X"00000001";

	when X"800009a8" => n_pc <= X"800009ac"; 
 if unsigned(reg8) >= unsigned(reg24) then n_pc <= X"800009b0"; end if;

	when X"800009ac" => n_pc <= X"800009b0"; 
 if signed(reg8) /= signed(reg13) then n_pc <= X"80000998"; end if;

	when X"800009b0" => n_pc <= X"800009b4"; 
 n_reg13 <= X"0000001f";

	when X"800009b4" => n_pc <= X"800009b8"; 
 n_reg12 <= X"00000030";

	when X"800009b8" => n_pc <= X"800009bc"; 
 if signed(reg14) = X"00000000" then n_pc <= X"800009c4"; end if;

	when X"800009bc" => n_pc <= X"800009c0"; 
 if unsigned(reg8) >= unsigned(reg26) then n_pc <= X"800009c4"; end if;

	when X"800009c0" => n_pc <= X"800009c4"; 
 if unsigned(reg13) >= unsigned(reg8) then n_pc <= X"80000a14"; end if;

	when X"800009c4" => n_pc <= X"800009c8"; 
 n_reg14 <= reg9 and X"00000010";

	when X"800009c8" => n_pc <= X"800009cc"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000a74"; end if;

	when X"800009cc" => n_pc <= X"800009d0"; 
 if signed(reg25) /= X"00000000" then n_pc <= X"80000a2c"; end if;

	when X"800009d0" => n_pc <= X"800009d4"; 
 if signed(reg8) = X"00000000" then n_pc <= X"80000a2c"; end if;

	when X"800009d4" => n_pc <= X"800009d8"; 
 if signed(reg24) = signed(reg8) then n_pc <= X"800009dc"; end if;

	when X"800009d8" => n_pc <= X"800009dc"; 
 if signed(reg8) /= signed(reg26) then n_pc <= X"80000a2c"; end if;

	when X"800009dc" => n_pc <= X"800009e0"; 
 n_reg14 <= reg8 + X"ffffffff";

	when X"800009e0" => n_pc <= X"800009e4"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000a28"; end if;

	when X"800009e4" => n_pc <= X"800009e8"; 
 n_reg13 <= X"00000010";

	when X"800009e8" => n_pc <= X"800009ec"; 
 n_reg8 <= reg8 + X"fffffffe";

	when X"800009ec" => n_pc <= X"800009f0"; 
 if signed(reg11) = signed(reg13) then n_pc <= X"80000a34"; end if;

	when X"800009f0" => n_pc <= X"800009f4"; 
 n_reg8 <= reg14;

	when X"800009f4" => n_pc <= X"800009f8"; 
 n_reg14 <= X"00000002";

	when X"800009f8" => n_pc <= X"800009fc"; 
 if signed(reg11) /= signed(reg14) then n_pc <= X"80000a58"; end if;

	when X"800009fc" => n_pc <= X"80000a00"; 
 n_reg14 <= X"0000001f";

	when X"80000a00" => n_pc <= X"80000a04"; 
 if unsigned(reg14) < unsigned(reg8) then n_pc <= X"80000a98"; end if;

	when X"80000a04" => n_pc <= X"80000a08"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000a08" => n_pc <= X"80000a0c"; 
 n_reg14 <= reg15 + reg8;

	when X"80000a0c" => n_pc <= X"80000a10"; 
 n_reg13 <= X"00000062";

	when X"80000a10" => 
 n_pc <= X"80000a50";

	when X"80000a14" => n_pc <= X"80000a18"; 
 n_reg15 <= reg2 + X"00000010";

	when X"80000a18" => n_pc <= X"80000a1c"; 
 n_reg10 <= reg15 + reg8;

	when X"80000a1c" => mem_width <= "00"; n_mem_addr <= reg10; n_mem_wdata <= reg12; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000A20";
 end if;
	when X"80000a20" => n_pc <= X"80000a24"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000a24" => 
 n_pc <= X"800009b8";

	when X"80000a28" => n_pc <= X"80000a2c"; 
 n_reg8 <= X"00000000";

	when X"80000a2c" => n_pc <= X"80000a30"; 
 n_reg14 <= X"00000010";

	when X"80000a30" => n_pc <= X"80000a34"; 
 if signed(reg11) /= signed(reg14) then n_pc <= X"800009f4"; end if;

	when X"80000a34" => n_pc <= X"80000a38"; 
 n_reg14 <= reg9 and X"00000020";

	when X"80000a38" => n_pc <= X"80000a3c"; 
 if signed(reg14) /= X"00000000" then n_pc <= X"80000ab0"; end if;

	when X"80000a3c" => n_pc <= X"80000a40"; 
 n_reg14 <= X"0000001f";

	when X"80000a40" => n_pc <= X"80000a44"; 
 if unsigned(reg14) < unsigned(reg8) then n_pc <= X"80000a98"; end if;

	when X"80000a44" => n_pc <= X"80000a48"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000a48" => n_pc <= X"80000a4c"; 
 n_reg14 <= reg15 + reg8;

	when X"80000a4c" => n_pc <= X"80000a50"; 
 n_reg13 <= X"00000078";

	when X"80000a50" => mem_width <= "00"; n_mem_addr <= reg14 + X"00000fe0"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000A54";
 end if;
	when X"80000a54" => n_pc <= X"80000a58"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000a58" => n_pc <= X"80000a5c"; 
 n_reg14 <= X"0000001f";

	when X"80000a5c" => n_pc <= X"80000a60"; 
 if unsigned(reg14) < unsigned(reg8) then n_pc <= X"80000a98"; end if;

	when X"80000a60" => n_pc <= X"80000a64"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000a64" => n_pc <= X"80000a68"; 
 n_reg14 <= reg15 + reg8;

	when X"80000a68" => n_pc <= X"80000a6c"; 
 n_reg13 <= X"00000030";

	when X"80000a6c" => mem_width <= "00"; n_mem_addr <= reg14 + X"00000fe0"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000A70";
 end if;
	when X"80000a70" => n_pc <= X"80000a74"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000a74" => n_pc <= X"80000a78"; 
 n_reg14 <= X"0000001f";

	when X"80000a78" => n_pc <= X"80000a7c"; 
 if unsigned(reg14) < unsigned(reg8) then n_pc <= X"80000a98"; end if;

	when X"80000a7c" => n_mem_addr <= reg2 + X"00000008"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000A80"; n_reg15 <= (others => '0');n_reg15(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000a80" => n_pc <= X"80000a84"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000ac8"; end if;

	when X"80000a84" => n_pc <= X"80000a88"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000a88" => n_pc <= X"80000a8c"; 
 n_reg14 <= reg15 + reg8;

	when X"80000a8c" => n_pc <= X"80000a90"; 
 n_reg13 <= X"0000002d";

	when X"80000a90" => mem_width <= "00"; n_mem_addr <= reg14 + X"00000fe0"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000A94";
 end if;
	when X"80000a94" => n_pc <= X"80000a98"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000a98" => n_pc <= X"80000a9c"; 
 n_reg9 <= reg9 and X"00000003";

	when X"80000a9c" => n_pc <= X"80000aa0"; 
 n_reg24 <= reg18;

	when X"80000aa0" => n_pc <= X"80000aa4"; 
 if signed(reg9) /= X"00000000" then n_pc <= X"80000b24"; end if;

	when X"80000aa4" => n_pc <= X"80000aa8"; 
 n_reg9 <= reg8;

	when X"80000aa8" => n_pc <= X"80000aac"; 
 n_reg23 <= reg18 - reg8;

	when X"80000aac" => 
 n_pc <= X"80000b0c";

	when X"80000ab0" => n_pc <= X"80000ab4"; 
 n_reg14 <= X"0000001f";

	when X"80000ab4" => n_pc <= X"80000ab8"; 
 if unsigned(reg14) < unsigned(reg8) then n_pc <= X"80000a98"; end if;

	when X"80000ab8" => n_pc <= X"80000abc"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000abc" => n_pc <= X"80000ac0"; 
 n_reg14 <= reg15 + reg8;

	when X"80000ac0" => n_pc <= X"80000ac4"; 
 n_reg13 <= X"00000058";

	when X"80000ac4" => 
 n_pc <= X"80000a50";

	when X"80000ac8" => n_pc <= X"80000acc"; 
 n_reg14 <= reg9 and X"00000004";

	when X"80000acc" => n_pc <= X"80000ad0"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000ae0"; end if;

	when X"80000ad0" => n_pc <= X"80000ad4"; 
 n_reg15 <= reg2 + X"00000030";

	when X"80000ad4" => n_pc <= X"80000ad8"; 
 n_reg14 <= reg15 + reg8;

	when X"80000ad8" => n_pc <= X"80000adc"; 
 n_reg13 <= X"0000002b";

	when X"80000adc" => 
 n_pc <= X"80000a90";

	when X"80000ae0" => n_pc <= X"80000ae4"; 
 n_reg14 <= reg9 and X"00000008";

	when X"80000ae4" => n_pc <= X"80000ae8"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000a98"; end if;

	when X"80000ae8" => n_pc <= X"80000aec"; 
 n_reg15 <= reg2 + X"00000030";
	when X"80000aec" => n_pc <= X"80000af0"; 
 n_reg14 <= reg15 + reg8;

	when X"80000af0" => n_pc <= X"80000af4"; 
 n_reg13 <= X"00000020";

	when X"80000af4" => 
 n_pc <= X"80000a90";

	when X"80000af8" => n_pc <= X"80000afc"; 
 n_reg13 <= reg22;

	when X"80000afc" => n_pc <= X"80000b00"; 
 n_reg11 <= reg21;

	when X"80000b00" => n_pc <= X"80000b04"; 
 n_reg10 <= X"00000020";

	when X"80000b04" => 
 n_reg1 <= X"80000B08"; n_pc <= reg20 + X"00000000";

	when X"80000b08" => n_pc <= X"80000b0c"; 
 n_reg9 <= reg9 + X"00000001";

	when X"80000b0c" => n_pc <= X"80000b10"; 
 n_reg12 <= reg23 + reg9;

	when X"80000b10" => n_pc <= X"80000b14"; 
 if unsigned(reg9) < unsigned(reg26) then n_pc <= X"80000af8"; end if;

	when X"80000b14" => n_pc <= X"80000b18"; 
 n_reg24 <= X"00000000";

	when X"80000b18" => n_pc <= X"80000b1c"; 
 if unsigned(reg26) < unsigned(reg8) then n_pc <= X"80000b20"; end if;

	when X"80000b1c" => n_pc <= X"80000b20"; 
 n_reg24 <= reg26 - reg8;

	when X"80000b20" => n_pc <= X"80000b24"; 
 n_reg24 <= reg24 + reg18;

	when X"80000b24" => n_pc <= X"80000b28"; 
 n_reg23 <= reg8;

	when X"80000b28" => n_pc <= X"80000b2c"; 
 n_reg9 <= reg8 + reg24;

	when X"80000b2c" => n_pc <= X"80000b30"; 
 n_reg12 <= reg9 - reg23;

	when X"80000b30" => n_pc <= X"80000b34"; 
 if signed(reg23) /= X"00000000" then n_pc <= X"80000b9c"; end if;

	when X"80000b34" => n_pc <= X"80000b38"; 
 if signed(reg19) = X"00000000" then n_pc <= X"80000b5c"; end if;

	when X"80000b38" => n_pc <= X"80000b3c"; 
 n_reg19 <= reg9 - reg18;

	when X"80000b3c" => n_pc <= X"80000b40"; 
 n_reg8 <= reg19;

	when X"80000b40" => n_pc <= X"80000b44"; 
 n_reg12 <= reg18 + reg8;

	when X"80000b44" => n_pc <= X"80000b48"; 
 if unsigned(reg8) < unsigned(reg26) then n_pc <= X"80000bbc"; end if;

	when X"80000b48" => n_pc <= X"80000b4c"; 
 n_reg12 <= X"00000000";

	when X"80000b4c" => n_pc <= X"80000b50"; 
 if unsigned(reg26) < unsigned(reg19) then n_pc <= X"80000b58"; end if;

	when X"80000b50" => n_pc <= X"80000b54"; 
 n_reg18 <= reg18 + reg26;

	when X"80000b54" => n_pc <= X"80000b58"; 
 n_reg12 <= reg18 - reg9;

	when X"80000b58" => n_pc <= X"80000b5c"; 
 n_reg9 <= reg9 + reg12;

	when X"80000b5c" => n_mem_addr <= reg2 + X"0000006c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B60"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b60" => n_mem_addr <= reg2 + X"00000068"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B64"; n_reg8 <= (others => '0');n_reg8(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b64" => n_mem_addr <= reg2 + X"00000060"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B68"; n_reg18 <= (others => '0');n_reg18(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b68" => n_mem_addr <= reg2 + X"0000005c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B6C"; n_reg19 <= (others => '0');n_reg19(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b6c" => n_mem_addr <= reg2 + X"00000058"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B70"; n_reg20 <= (others => '0');n_reg20(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b70" => n_mem_addr <= reg2 + X"00000054"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B74"; n_reg21 <= (others => '0');n_reg21(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b74" => n_mem_addr <= reg2 + X"00000050"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B78"; n_reg22 <= (others => '0');n_reg22(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b78" => n_mem_addr <= reg2 + X"0000004c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B7C"; n_reg23 <= (others => '0');n_reg23(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b7c" => n_mem_addr <= reg2 + X"00000048"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B80"; n_reg24 <= (others => '0');n_reg24(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b80" => n_mem_addr <= reg2 + X"00000044"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B84"; n_reg25 <= (others => '0');n_reg25(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b84" => n_mem_addr <= reg2 + X"00000040"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B88"; n_reg26 <= (others => '0');n_reg26(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b88" => n_mem_addr <= reg2 + X"0000003c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B8C"; n_reg27 <= (others => '0');n_reg27(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b8c" => n_pc <= X"80000b90"; 
 n_reg10 <= reg9;

	when X"80000b90" => n_mem_addr <= reg2 + X"00000064"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000B94"; n_reg9 <= (others => '0');n_reg9(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000b94" => n_pc <= X"80000b98"; 
 n_reg2 <= reg2 + X"00000070";

	when X"80000b98" => 
 n_pc <= reg1;

	when X"80000b9c" => n_pc <= X"80000ba0"; 
 n_reg23 <= reg23 + X"ffffffff";

	when X"80000ba0" => n_pc <= X"80000ba4"; 
 n_reg15 <= reg2 + X"00000010";

	when X"80000ba4" => n_pc <= X"80000ba8"; 
 n_reg14 <= reg15 + reg23;

	when X"80000ba8" => n_mem_addr <= reg14; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000BAC"; n_reg10 <= (others => '0');n_reg10(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000bac" => n_pc <= X"80000bb0"; 
 n_reg13 <= reg22;

	when X"80000bb0" => n_pc <= X"80000bb4"; 
 n_reg11 <= reg21;

	when X"80000bb4" => 
 n_reg1 <= X"80000BB8"; n_pc <= reg20 + X"00000000";

	when X"80000bb8" => 
 n_pc <= X"80000b28";

	when X"80000bbc" => n_pc <= X"80000bc0"; 
 n_reg13 <= reg22;

	when X"80000bc0" => n_pc <= X"80000bc4"; 
 n_reg11 <= reg21;

	when X"80000bc4" => n_pc <= X"80000bc8"; 
 n_reg10 <= X"00000020";

	when X"80000bc8" => 
 n_reg1 <= X"80000BCC"; n_pc <= reg20 + X"00000000";

	when X"80000bcc" => n_pc <= X"80000bd0"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80000bd0" => 
 n_pc <= X"80000b40";

	when X"80000bd4" => n_pc <= X"80000bd8"; 
 if signed(reg10) = X"00000000" then n_pc <= X"80000bdc"; end if;

	when X"80000bd8" => 
 n_pc <= X"80000838";

	when X"80000bdc" => 
 n_pc <= reg1;

	when X"80000be0" => n_pc <= X"80000be4"; 
 if signed(reg10) = X"00000000" then n_pc <= X"80000bf0"; end if;

	when X"80000be4" => n_mem_addr <= reg11; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000BE8"; n_reg6 <= (others => '0');n_reg6(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000be8" => n_mem_addr <= reg11 + X"00000004"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000BEC"; n_reg11 <= (others => '0');n_reg11(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000bec" => 
 n_pc <= reg6;

	when X"80000bf0" => 
 n_pc <= reg1;

	when X"80000bf4" => n_pc <= X"80000bf8"; 
 n_reg2 <= reg2 + X"ffffffa0";

	when X"80000bf8" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000054"; n_mem_wdata <= reg9; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000BFC";
 end if;
	when X"80000bfc" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000050"; n_mem_wdata <= reg18; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C00";
 end if;
	when X"80000c00" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000004c"; n_mem_wdata <= reg19; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C04";
 end if;
	when X"80000c04" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000048"; n_mem_wdata <= reg20; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C08";
 end if;
	when X"80000c08" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg23; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C0C";
 end if;
	when X"80000c0c" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000005c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C10";
 end if;
	when X"80000c10" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000058"; n_mem_wdata <= reg8; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C14";
 end if;
	when X"80000c14" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000044"; n_mem_wdata <= reg21; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C18";
 end if;
	when X"80000c18" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000040"; n_mem_wdata <= reg22; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C1C";
 end if;
	when X"80000c1c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000038"; n_mem_wdata <= reg24; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C20";
 end if;
	when X"80000c20" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000034"; n_mem_wdata <= reg25; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C24";
 end if;
	when X"80000c24" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000030"; n_mem_wdata <= reg26; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000C28";
 end if;
	when X"80000c28" => 
		mem_width <= "10"; 
		n_mem_addr <= reg2 + X"0000002c"; 
		n_mem_wdata <= reg27; 
		mem_we <= '1'; 
		if mem_wack = '1' then
			n_pc <= X"80000C2C";
		end if;
	when X"80000c2c" => 
	n_pc <= X"80000c30"; 
 	n_reg20 <= reg11;

	when X"80000c30" => n_pc <= X"80000c34"; 
 n_reg19 <= reg12;

	when X"80000c34" => n_pc <= X"80000c38"; 
 n_reg9 <= reg13;

	when X"80000c38" => n_pc <= X"80000c3c"; 
 n_reg23 <= reg14;
	when X"80000c3c" => n_pc <= X"80000c40"; 
 n_reg18 <= reg10;

	when X"80000c40" => n_pc <= X"80000c44"; 
 if signed(reg11) /= X"00000000" then n_pc <= X"80000c4c"; end if;

	when X"80000c44" => n_pc <= X"80000c48"; 
 n_reg18 <= X"80001000";

	when X"80000c48" => n_pc <= X"80000c4c"; 
 n_reg18 <= reg18 + X"fffff870";

	when X"80000c4c" => 
		n_pc <= X"80000c50"; 
		n_reg21 <= X"00010000";

	when X"80000c50" => n_pc <= X"80000c54"; 
 n_reg22 <= X"80000000";

	when X"80000c54" => n_pc <= X"80000c58"; 
 n_reg27 <= X"00000000";

	when X"80000c58" => n_pc <= X"80000c5c"; 
 n_reg21 <= reg21 + X"ffffffff";

	when X"80000c5c" => n_pc <= X"80000c60"; 
 n_reg22 <= reg22 + X"00000010";

	when X"80000c60" => 
 n_pc <= X"80001074";

	when X"80000c64" => n_pc <= X"80000c68"; 
 n_reg15 <= X"00000025";

	when X"80000c68" => n_pc <= X"80000c6c"; 
 n_reg9 <= reg9 + X"00000001";

	when X"80000c6c" => n_pc <= X"80000c70"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80000c84"; end if;

	when X"80000c70" => n_pc <= X"80000c74"; 
 n_reg8 <= reg27 + X"00000001";

	when X"80000c74" => n_pc <= X"80000c78"; 
 n_reg13 <= reg19;

	when X"80000c78" => n_pc <= X"80000c7c"; 
 n_reg12 <= reg27;

	when X"80000c7c" => n_pc <= X"80000c80"; 
 n_reg11 <= reg20;

	when X"80000c80" => 
 n_pc <= X"8000125c";

	when X"80000c84" => n_pc <= X"80000c88"; 
 n_reg6 <= X"00000000";

	when X"80000c88" => n_pc <= X"80000c8c"; 
 n_reg14 <= X"0000002b";

	when X"80000c8c" => n_pc <= X"80000c90"; 
 n_reg12 <= X"00000020";

	when X"80000c90" => n_pc <= X"80000c94"; 
 n_reg11 <= X"00000023";

	when X"80000c94" => 
 n_pc <= X"80000cb0";

	when X"80000c98" => n_pc <= X"80000c9c"; 
 n_reg10 <= X"0000002d";

	when X"80000c9c" => n_pc <= X"80000ca0"; 
 if signed(reg15) = signed(reg10) then n_pc <= X"80000ce4"; end if;

	when X"80000ca0" => n_pc <= X"80000ca4"; 
 n_reg10 <= X"00000030";

	when X"80000ca4" => n_pc <= X"80000ca8"; 
 if signed(reg15) /= signed(reg10) then n_pc <= X"80000cc8"; end if;

	when X"80000ca8" => n_pc <= X"80000cac"; 
 n_reg6 <= reg6 or X"00000001";

	when X"80000cac" => n_pc <= X"80000cb0"; 
 n_reg9 <= reg13;

	when X"80000cb0" => n_mem_addr <= reg9; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000CB4"; n_reg15 <= (others => '0');n_reg15(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000cb4" => n_pc <= X"80000cb8"; 
 n_reg13 <= reg9 + X"00000001";

	when X"80000cb8" => n_pc <= X"80000cbc"; 
 if signed(reg15) = signed(reg14) then n_pc <= X"80000cec"; end if;

	when X"80000cbc" => n_pc <= X"80000cc0"; 
 if unsigned(reg14) < unsigned(reg15) then n_pc <= X"80000c98"; end if;

	when X"80000cc0" => n_pc <= X"80000cc4"; 
 if signed(reg15) = signed(reg12) then n_pc <= X"80000cf4"; end if;

	when X"80000cc4" => n_pc <= X"80000cc8"; 
 if signed(reg15) = signed(reg11) then n_pc <= X"80000cfc"; end if;

	when X"80000cc8" => n_pc <= X"80000ccc"; 
 n_reg14 <= reg15 + X"ffffffd0";

	when X"80000ccc" => n_pc <= X"80000cd0"; 
 n_reg14 <= reg14 and X"000000ff";

	when X"80000cd0" => n_pc <= X"80000cd4"; 
 n_reg12 <= X"00000009";

	when X"80000cd4" => n_pc <= X"80000cd8"; 
 if unsigned(reg12) < unsigned(reg14) then n_pc <= X"80000d64"; end if;

	when X"80000cd8" => n_pc <= X"80000cdc"; 
 n_reg24 <= X"00000000";

	when X"80000cdc" => n_pc <= X"80000ce0"; 
 n_reg13 <= X"00000009";

	when X"80000ce0" => 
 n_pc <= X"80000d1c";

	when X"80000ce4" => n_pc <= X"80000ce8"; 
 n_reg6 <= reg6 or X"00000002";

	when X"80000ce8" => 
 n_pc <= X"80000cac";

	when X"80000cec" => n_pc <= X"80000cf0"; 
 n_reg6 <= reg6 or X"00000004";

	when X"80000cf0" => 
 n_pc <= X"80000cac";

	when X"80000cf4" => n_pc <= X"80000cf8"; 
 n_reg6 <= reg6 or X"00000008";

	when X"80000cf8" => 
 n_pc <= X"80000cac";

	when X"80000cfc" => n_pc <= X"80000d00"; 
 n_reg6 <= reg6 or X"00000010";

	when X"80000d00" => 
 n_pc <= X"80000cac";

	when X"80000d04" => n_pc <= X"80000d08"; 
 n_reg15 <= (others => '0'); n_reg15(31 downto 2) <= reg24(29 downto 0);

	when X"80000d08" => n_pc <= X"80000d0c"; 
 n_reg28 <= reg15 + reg24;

	when X"80000d0c" => n_pc <= X"80000d10"; 
 n_reg28 <= (others => '0'); n_reg28(31 downto 1) <= reg28(30 downto 0);

	when X"80000d10" => n_pc <= X"80000d14"; 
 n_reg28 <= reg28 + X"ffffffd0";

	when X"80000d14" => n_pc <= X"80000d18"; 
 n_reg24 <= reg14 + reg28;

	when X"80000d18" => n_pc <= X"80000d1c"; 
 n_reg9 <= reg12;

	when X"80000d1c" => n_mem_addr <= reg9; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000D20"; n_reg14 <= (others => '0');n_reg14(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000d20" => n_pc <= X"80000d24"; 
 n_reg12 <= reg9 + X"00000001";

	when X"80000d24" => n_pc <= X"80000d28"; 
 n_reg15 <= reg14 + X"ffffffd0";

	when X"80000d28" => n_pc <= X"80000d2c"; 
 n_reg15 <= reg15 and X"000000ff";

	when X"80000d2c" => n_pc <= X"80000d30"; 
 if unsigned(reg13) >= unsigned(reg15) then n_pc <= X"80000d04"; end if;

	when X"80000d30" => n_mem_addr <= reg9; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000D34"; n_reg14 <= (others => '0');n_reg14(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000d34" => n_pc <= X"80000d38"; 
 n_reg15 <= X"0000002e";

	when X"80000d38" => n_pc <= X"80000d3c"; 
 n_reg17 <= X"00000000";

	when X"80000d3c" => n_pc <= X"80000d40"; 
 if signed(reg14) /= signed(reg15) then n_pc <= X"80000de4"; end if;

	when X"80000d40" => n_mem_addr <= reg9 + X"00000001"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000D44"; n_reg13 <= (others => '0');n_reg13(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000d44" => n_pc <= X"80000d48"; 
 n_reg12 <= X"00000009";

	when X"80000d48" => n_pc <= X"80000d4c"; 
 n_reg15 <= reg9 + X"00000001";

	when X"80000d4c" => n_pc <= X"80000d50"; 
 n_reg14 <= reg13 + X"ffffffd0";

	when X"80000d50" => n_pc <= X"80000d54"; 
 n_reg14 <= reg14 and X"000000ff";

	when X"80000d54" => n_pc <= X"80000d58"; 
 n_reg6 <= reg6 or X"00000400";

	when X"80000d58" => n_pc <= X"80000d5c";
 if unsigned(reg12) < unsigned(reg14) then n_pc <= X"80000dc4"; end if;

	when X"80000d5c" => n_pc <= X"80000d60"; 
 n_reg12 <= X"00000009";

	when X"80000d60" => 
 n_pc <= X"80000da8";

	when X"80000d64" => n_pc <= X"80000d68"; 
 n_reg14 <= X"0000002a";

	when X"80000d68" => n_pc <= X"80000d6c"; 
 n_reg24 <= X"00000000";

	when X"80000d6c" => n_pc <= X"80000d70"; 
 if signed(reg15) /= signed(reg14) then n_pc <= X"80000d30"; end if;

	when X"80000d70" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000D74"; n_reg24 <= (others => '0');n_reg24(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000d74" => n_pc <= X"80000d78"; 
 n_reg15 <= reg23 + X"00000004";

	when X"80000d78" => n_pc <= X"80000d7c";
 if signed(reg24) >= X"00000000" then n_pc <= X"80000d84"; end if;

	when X"80000d7c" => n_pc <= X"80000d80"; 
 n_reg6 <= reg6 or X"00000002";

	when X"80000d80" => n_pc <= X"80000d84"; 
 n_reg24 <= X"00000000" - reg24;

	when X"80000d84" => n_pc <= X"80000d88"; 
 n_reg23 <= reg15;

	when X"80000d88" => n_pc <= X"80000d8c"; 
 n_reg9 <= reg13;

	when X"80000d8c" => 
 n_pc <= X"80000d30";

	when X"80000d90" => n_pc <= X"80000d94"; 
 n_reg15 <= (others => '0'); n_reg15(31 downto 2) <= reg17(29 downto 0);

	when X"80000d94" => n_pc <= X"80000d98"; 
 n_reg17 <= reg15 + reg17;

	when X"80000d98" => n_pc <= X"80000d9c"; 
 n_reg17 <= (others => '0'); n_reg17(31 downto 1) <= reg17(30 downto 0);

	when X"80000d9c" => n_pc <= X"80000da0"; 
 n_reg17 <= reg17 + X"ffffffd0";

	when X"80000da0" => n_pc <= X"80000da4"; 
 n_reg17 <= reg13 + reg17;

	when X"80000da4" => n_pc <= X"80000da8"; 
 n_reg15 <= reg11;

	when X"80000da8" => n_mem_addr <= reg15; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000DAC"; n_reg13 <= (others => '0');n_reg13(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000dac" => n_pc <= X"80000db0"; 
 n_reg11 <= reg15 + X"00000001";

	when X"80000db0" => n_pc <= X"80000db4"; 
 n_reg14 <= reg13 + X"ffffffd0";

	when X"80000db4" => n_pc <= X"80000db8"; 
 n_reg14 <= reg14 and X"000000ff";

	when X"80000db8" => n_pc <= X"80000dbc"; 
 if unsigned(reg12) >= unsigned(reg14) then n_pc <= X"80000d90"; end if;

	when X"80000dbc" => n_pc <= X"80000dc0"; 
 n_reg9 <= reg15;

	when X"80000dc0" => 
 n_pc <= X"80000de4";

	when X"80000dc4" => n_pc <= X"80000dc8"; 
 n_reg14 <= X"0000002a";

	when X"80000dc8" => n_pc <= X"80000dcc"; 
 if signed(reg13) /= signed(reg14) then n_pc <= X"80000dbc"; end if;

	when X"80000dcc" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000DD0"; n_reg17 <= (others => '0');n_reg17(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000dd0" => n_pc <= X"80000dd4"; 
 n_reg15 <= reg23 + X"00000004";

	when X"80000dd4" => n_pc <= X"80000dd8"; 
 if signed(reg17) >= X"00000000" then n_pc <= X"80000ddc"; end if;

	when X"80000dd8" => n_pc <= X"80000ddc"; 
 n_reg17 <= X"00000000";

	when X"80000ddc" => n_pc <= X"80000de0"; 
 n_reg9 <= reg9 + X"00000002";

	when X"80000de0" => n_pc <= X"80000de4"; 
 n_reg23 <= reg15;

	when X"80000de4" => n_mem_addr <= reg9; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000DE8"; n_reg15 <= (others => '0');n_reg15(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000de8" => n_pc <= X"80000dec"; 
 n_reg13 <= X"0000006c";

	when X"80000dec" => n_pc <= X"80000df0"; 
 n_reg14 <= reg9 + X"00000001";

	when X"80000df0" => n_pc <= X"80000df4"; 
 if signed(reg15) = signed(reg13) then n_pc <= X"80000e58"; end if;

	when X"80000df4" => n_pc <= X"80000df8"; 
 if unsigned(reg13) < unsigned(reg15) then n_pc <= X"80000e40"; end if;

	when X"80000df8" => n_pc <= X"80000dfc"; 
 n_reg13 <= X"00000068";

	when X"80000dfc" => n_pc <= X"80000e00"; 
 if signed(reg15) = signed(reg13) then n_pc <= X"80000e6c"; end if;

	when X"80000e00" => n_pc <= X"80000e04"; 
 n_reg13 <= X"0000006a";

	when X"80000e04" => n_pc <= X"80000e08"; 
 if signed(reg15) = signed(reg13) then n_pc <= X"80000e84"; end if;

	when X"80000e08" => n_pc <= X"80000e0c"; 
 n_reg14 <= reg9;

	when X"80000e0c" => n_mem_addr <= reg14; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000E10"; n_reg10 <= (others => '0');n_reg10(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000e10" => n_pc <= X"80000e14"; 
 n_reg15 <= X"00000078";

	when X"80000e14" => n_pc <= X"80000e18"; 
 n_reg9 <= reg14 + X"00000001";

	when X"80000e18" => n_pc <= X"80000e1c"; 
 if unsigned(reg15) < unsigned(reg10) then n_pc <= X"80000c70"; end if;

	when X"80000e1c" => n_pc <= X"80000e20"; 
 n_reg15 <= X"00000061";

	when X"80000e20" => n_pc <= X"80000e24"; 
 if unsigned(reg15) < unsigned(reg10) then n_pc <= X"80000e8c"; end if;

	when X"80000e24" => n_pc <= X"80000e28"; 
 n_reg15 <= X"00000025";

	when X"80000e28" => n_pc <= X"80000e2c"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80001248"; end if;

	when X"80000e2c" => n_pc <= X"80000e30"; 
 n_reg15 <= X"00000058";

	when X"80000e30" => n_pc <= X"80000e34"; 
 if signed(reg10) /= signed(reg15) then n_pc <= X"80000c70"; end if;

	when X"80000e34" => n_pc <= X"80000e38"; 
 n_reg6 <= reg6 or X"00000020";

	when X"80000e38" => n_pc <= X"80000e3c"; 
 n_reg16 <= X"00000010";

	when X"80000e3c" => 
 n_pc <= X"80000edc";

	when X"80000e40" => n_pc <= X"80000e44"; 
 n_reg13 <= X"00000074";

	when X"80000e44" => n_pc <= X"80000e48"; 
 if signed(reg15) = signed(reg13) then n_pc <= X"80000e50"; end if;

	when X"80000e48" => n_pc <= X"80000e4c"; 
 n_reg13 <= X"0000007a";

	when X"80000e4c" => n_pc <= X"80000e50"; 
 if signed(reg15) /= signed(reg13) then n_pc <= X"80000e08"; end if;

	when X"80000e50" => n_pc <= X"80000e54"; 
 n_reg6 <= reg6 or X"00000100";

	when X"80000e54" => 
 n_pc <= X"80000e0c";

	when X"80000e58" => n_mem_addr <= reg9 + X"00000001"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000E5C"; n_reg13 <= (others => '0');n_reg13(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000e5c" => n_pc <= X"80000e60"; 
 if signed(reg13) /= signed(reg15) then n_pc <= X"80000e50"; end if;

	when X"80000e60" => n_pc <= X"80000e64"; 
 n_reg6 <= reg6 or X"00000300";

	when X"80000e64" => n_pc <= X"80000e68"; 
 n_reg14 <= reg9 + X"00000002";

	when X"80000e68" => 
 n_pc <= X"80000e0c";

	when X"80000e6c" => n_mem_addr <= reg9 + X"00000001"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000E70"; n_reg13 <= (others => '0');n_reg13(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80000e70" => n_pc <= X"80000e74"; 
 if signed(reg13) = signed(reg15) then n_pc <= X"80000e7c"; end if;

	when X"80000e74" => n_pc <= X"80000e78"; 
 n_reg6 <= reg6 or X"00000080";

	when X"80000e78" => 
 n_pc <= X"80000e0c";

	when X"80000e7c" => n_pc <= X"80000e80"; 
 n_reg6 <= reg6 or X"000000c0";

	when X"80000e80" => 
 n_pc <= X"80000e64";

	when X"80000e84" => n_pc <= X"80000e88"; 
 n_reg6 <= reg6 or X"00000200";

	when X"80000e88" => 
 n_pc <= X"80000e0c";

	when X"80000e8c" => n_pc <= X"80000e90"; 
 n_reg15 <= reg10 + X"ffffff9e";

	when X"80000e90" => n_pc <= X"80000e94"; 
 n_reg15 <= reg15 and X"000000ff";

	when X"80000e94" => n_pc <= X"80000e98"; 
 n_reg14 <= X"00000016";

	when X"80000e98" => n_pc <= X"80000e9c"; 
 if unsigned(reg14) < unsigned(reg15) then n_pc <= X"80000c70"; end if;

	when X"80000e9c" => n_pc <= X"80000ea0"; 
 n_reg15 <= (others => '0'); n_reg15(31 downto 2) <= reg15(29 downto 0);

	when X"80000ea0" => n_pc <= X"80000ea4"; 
 n_reg15 <= reg15 + reg22;

	when X"80000ea4" => n_mem_addr <= reg15; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000EA8"; n_reg15 <= (others => '0');n_reg15(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000ea8" => 
 n_pc <= reg15;

	when X"80000eac" => n_pc <= X"80000eb0"; 
 n_reg15 <= X"00000078";

	when X"80000eb0" => n_pc <= X"80000eb4"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80000e38"; end if;

	when X"80000eb4" => n_pc <= X"80000eb8"; 
 n_reg15 <= X"0000006f";

	when X"80000eb8" => n_pc <= X"80000ebc"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80001268"; end if;

	when X"80000ebc" => n_pc <= X"80000ec0"; 
 n_reg15 <= X"00000062";

	when X"80000ec0" => n_pc <= X"80000ec4"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80001270"; end if;

	when X"80000ec4" => n_pc <= X"80000ec8"; 
 n_reg15 <= X"00000069";

	when X"80000ec8" => n_pc <= X"80000ecc"; 
 n_reg6 <= reg6 and X"ffffffef";

	when X"80000ecc" => n_pc <= X"80000ed0"; 
 n_reg16 <= X"0000000a";

	when X"80000ed0" => n_pc <= X"80000ed4"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80000ee0"; end if;

	when X"80000ed4" => n_pc <= X"80000ed8"; 
 n_reg15 <= X"00000064";

	when X"80000ed8" => n_pc <= X"80000edc"; 
 if signed(reg10) = signed(reg15) then n_pc <= X"80000ee0"; end if;

	when X"80000edc" => n_pc <= X"80000ee0"; 
 n_reg6 <= reg6 and X"fffffff3";

	when X"80000ee0" => n_pc <= X"80000ee4"; 
 n_reg15 <= reg6 and X"00000400";

	when X"80000ee4" => n_pc <= X"80000ee8"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000eec"; end if;

	when X"80000ee8" => n_pc <= X"80000eec"; 
 n_reg6 <= reg6 and X"fffffffe";

	when X"80000eec" => n_pc <= X"80000ef0"; 
 n_reg14 <= X"00000069";

	when X"80000ef0" => n_pc <= X"80000ef4"; 
 n_reg15 <= reg6 and X"00000200";

	when X"80000ef4" => n_pc <= X"80000ef8"; 
 if signed(reg10) = signed(reg14) then n_pc <= X"80000f00"; end if;

	when X"80000ef8" => n_pc <= X"80000efc"; 
 n_reg14 <= X"00000064";

	when X"80000efc" => n_pc <= X"80000f00"; 
 if signed(reg10) /= signed(reg14) then n_pc <= X"80000f74"; end if;

	when X"80000f00" => n_pc <= X"80000f04"; 
 if signed(reg15) /= X"00000000" then n_pc <= X"80001074"; end if;

	when X"80000f04" => n_pc <= X"80000f08"; 
 n_reg15 <= reg6 and X"00000100";

	when X"80000f08" => n_pc <= X"80000f0c"; 
 n_reg8 <= reg23 + X"00000004";

	when X"80000f0c" => n_pc <= X"80000f10"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000f4c"; end if;

	when X"80000f10" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000F14"; n_reg15 <= (others => '0');n_reg15(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000f14" => n_pc <= X"80000f18"; 
 n_reg15 <= (others => reg14(31)); n_reg14(0 downto 0) <= reg15(31 downto 31);

	when X"80000f18" => n_pc <= X"80000f1c"; 
 n_reg13 <= reg14 xor reg15;

	when X"80000f1c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000004"; n_mem_wdata <= reg6; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000F20";
 end if;
	when X"80000f20" => mem_width <= "10"; n_mem_addr <= reg2; n_mem_wdata <= reg24; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000F24";
 end if;
	when X"80000f24" => n_pc <= X"80000f28"; 
 n_reg15 <= (others => '0'); n_reg15(0 downto 0) <= reg15(31 downto 31);

	when X"80000f28" => n_pc <= X"80000f2c"; 
 n_reg14 <= reg13 - reg14;

	when X"80000f2c" => n_pc <= X"80000f30"; 
 n_reg12 <= reg27;

	when X"80000f30" => n_pc <= X"80000f34"; 
 n_reg13 <= reg19;

	when X"80000f34" => n_pc <= X"80000f38"; 
 n_reg11 <= reg20;

	when X"80000f38" => n_pc <= X"80000f3c"; 
 n_reg10 <= reg18;

	when X"80000f3c" => 
 n_reg1 <= X"80000F40"; n_pc <= X"80000874";

	when X"80000f40" => n_pc <= X"80000f44"; 
 n_reg27 <= reg10;

	when X"80000f44" => n_pc <= X"80000f48"; 
 n_reg23 <= reg8;

	when X"80000f48" => 
 n_pc <= X"80001074";

	when X"80000f4c" => n_pc <= X"80000f50"; 
 n_reg14 <= reg6 and X"00000040";

	when X"80000f50" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000F54"; n_reg15 <= (others => '0');n_reg15(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000f54" => n_pc <= X"80000f58"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000f60"; end if;

	when X"80000f58" => n_pc <= X"80000f5c"; 
 n_reg15 <= reg15 and X"000000ff";

	when X"80000f5c" => 
 n_pc <= X"80000f14";

	when X"80000f60" => n_pc <= X"80000f64"; 
 n_reg14 <= reg6 and X"00000080";

	when X"80000f64" => n_pc <= X"80000f68"; 
 if signed(reg14) = X"00000000" then n_pc <= X"80000f14"; end if;

	when X"80000f68" => n_pc <= X"80000f6c"; 
 n_reg15 <= (others => '0'); n_reg15(31 downto 16) <= reg15(15 downto 0);

	when X"80000f6c" => n_pc <= X"80000f70"; 
 n_reg15 <= (others => reg15(31)); n_reg15(15 downto 0) <= reg15(31 downto 16);

	when X"80000f70" => 
 n_pc <= X"80000f14";

	when X"80000f74" => n_pc <= X"80000f78"; 
 if signed(reg15) /= X"00000000" then n_pc <= X"80001074"; end if;

	when X"80000f78" => n_pc <= X"80000f7c"; 
 n_reg15 <= reg6 and X"00000100";

	when X"80000f7c" => n_pc <= X"80000f80"; 
 n_reg8 <= reg23 + X"00000004";

	when X"80000f80" => n_pc <= X"80000f84"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000f98"; end if;

	when X"80000f84" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000F88"; n_reg14 <= (others => '0');n_reg14(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000f88" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000004"; n_mem_wdata <= reg6; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000F8C";
 end if;
	when X"80000f8c" => mem_width <= "10"; n_mem_addr <= reg2; n_mem_wdata <= reg24; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80000F90";
 end if;
	when X"80000f90" => n_pc <= X"80000f94"; 
 n_reg15 <= X"00000000";

	when X"80000f94" => 
 n_pc <= X"80000f2c";

	when X"80000f98" => n_pc <= X"80000f9c"; 
 n_reg15 <= reg6 and X"00000040";

	when X"80000f9c" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80000FA0"; n_reg14 <= (others => '0');n_reg14(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80000fa0" => n_pc <= X"80000fa4"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000fac"; end if;

	when X"80000fa4" => n_pc <= X"80000fa8"; 
 n_reg14 <= reg14 and X"000000ff";

	when X"80000fa8" => 
 n_pc <= X"80000f88";

	when X"80000fac" => n_pc <= X"80000fb0"; 
 n_reg15 <= reg6 and X"00000080";

	when X"80000fb0" => n_pc <= X"80000fb4"; 
 if signed(reg15) = X"00000000" then n_pc <= X"80000f88"; end if;

	when X"80000fb4" => n_pc <= X"80000fb8"; 
 n_reg14 <= reg14 and reg21;

	when X"80000fb8" => 
 n_pc <= X"80000f88";

	when X"80000fbc" => n_pc <= X"80000fc0"; 
 n_reg8 <= reg6 and X"00000002";

	when X"80000fc0" => n_pc <= X"80000fc4"; 
 n_reg26 <= X"00000001";

	when X"80000fc4" => n_pc <= X"80000fc8"; 
 if signed(reg8) /= X"00000000" then n_pc <= X"8000100c"; end if;

	when X"80000fc8" => n_pc <= X"80000fcc"; 
 n_reg26 <= X"00000000";

	when X"80000fcc" => 
 n_pc <= X"80000fe0";

	when X"80000fd0" => n_pc <= X"80000fd4"; 
 n_reg13 <= reg19;

	when X"80000fd4" => n_pc <= X"80000fd8"; 
 n_reg11 <= reg20;

	when X"80000fd8" => n_pc <= X"80000fdc"; 
 n_reg10 <= X"00000020";

	when X"80000fdc" => 
 n_reg1 <= X"80000FE0"; n_pc <= reg18 + X"00000000";

	when X"80000fe0" => n_pc <= X"80000fe4"; 
 n_reg12 <= reg26 + reg27;

	when X"80000fe4" => n_pc <= X"80000fe8"; 
 n_reg26 <= reg26 + X"00000001";

	when X"80000fe8" => n_pc <= X"80000fec"; 
 if unsigned(reg26) < unsigned(reg24) then n_pc <= X"80000fd0"; end if;

	when X"80000fec" => n_pc <= X"80000ff0"; 
 n_reg15 <= X"00000000";

	when X"80000ff0" => n_pc <= X"80000ff4"; 
 if signed(reg24) = X"00000000" then n_pc <= X"80000ff8"; end if;

	when X"80000ff4" => n_pc <= X"80000ff8"; 
 n_reg15 <= reg24 + X"ffffffff";

	when X"80000ff8" => n_pc <= X"80000ffc"; 
 n_reg27 <= reg27 + reg15;

	when X"80000ffc" => n_pc <= X"80001000"; 
 n_reg15 <= X"00000002";

	when X"80001000" => n_pc <= X"80001004"; 
 if signed(reg24) = X"00000000" then n_pc <= X"80001008"; end if;

	when X"80001004" => n_pc <= X"80001008"; 
 n_reg15 <= reg24 + X"00000001";

	when X"80001008" => n_pc <= X"8000100c"; 
 n_reg26 <= reg15;

	when X"8000100c" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001010"; n_reg10 <= (others => '0');n_reg10(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80001010" => n_pc <= X"80001014"; 
 n_reg15 <= reg23 + X"00000004";

	when X"80001014" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000010"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001018";
 end if;
	when X"80001018" => n_pc <= X"8000101c"; 
 n_reg13 <= reg19;

	when X"8000101c" => n_pc <= X"80001020"; 
 n_reg12 <= reg27;

	when X"80001020" => n_pc <= X"80001024"; 
 n_reg11 <= reg20;

	when X"80001024" => n_pc <= X"80001028"; 
 n_reg25 <= reg27 + X"00000001";

	when X"80001028" => 
 n_reg1 <= X"8000102C"; n_pc <= reg18 + X"00000000";

	when X"8000102c" => n_pc <= X"80001030"; 
 if signed(reg8) = X"00000000" then n_pc <= X"8000106c"; end if;

	when X"80001030" => n_pc <= X"80001034"; 
 n_reg8 <= reg26;

	when X"80001034" => n_pc <= X"80001038"; 
 n_reg12 <= reg25;

	when X"80001038" => 
 n_pc <= X"80001058";

	when X"8000103c" => n_pc <= X"80001040"; 
 n_reg13 <= reg19;

	when X"80001040" => n_pc <= X"80001044"; 
 n_reg11 <= reg20;

	when X"80001044" => n_pc <= X"80001048"; 
 n_reg10 <= X"00000020";

	when X"80001048" => n_pc <= X"8000104c"; 
 n_reg23 <= reg12 + X"00000001";

	when X"8000104c" => 
 n_reg1 <= X"80001050"; n_pc <= reg18 + X"00000000";

	when X"80001050" => n_pc <= X"80001054"; 
 n_reg8 <= reg8 + X"00000001";

	when X"80001054" => n_pc <= X"80001058"; 
 n_reg12 <= reg23;

	when X"80001058" => n_pc <= X"8000105c"; 
 if unsigned(reg8) < unsigned(reg24) then n_pc <= X"8000103c"; end if;

	when X"8000105c" => n_pc <= X"80001060"; 
 n_reg13 <= X"00000000";

	when X"80001060" => n_pc <= X"80001064"; 
 if unsigned(reg24) < unsigned(reg26) then n_pc <= X"80001068"; end if;

	when X"80001064" => n_pc <= X"80001068"; 
 n_reg13 <= reg24 - reg26;

	when X"80001068" => n_pc <= X"8000106c"; 
 n_reg25 <= reg25 + reg13;

	when X"8000106c" => n_mem_addr <= reg2 + X"00000010"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001070"; n_reg23 <= (others => '0');n_reg23(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001070" => n_pc <= X"80001074"; 
 n_reg27 <= reg25;

	when X"80001074" => n_mem_addr <= reg9; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001078"; n_reg10 <= (others => '0');n_reg10(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"80001078" => n_pc <= X"8000107c"; 
 if signed(reg10) /= X"00000000" then n_pc <= X"80000c64"; end if;

	when X"8000107c" => n_pc <= X"80001080"; 
 n_reg12 <= reg27;

	when X"80001080" => n_pc <= X"80001084"; 
 if unsigned(reg27) < unsigned(reg19) then n_pc <= X"80001088"; end if;

	when X"80001084" => n_pc <= X"80001088"; 
 n_reg12 <= reg19 + X"ffffffff";

	when X"80001088" => n_pc <= X"8000108c"; 
 n_reg13 <= reg19;

	when X"8000108c" => n_pc <= X"80001090"; 
 n_reg11 <= reg20;

	when X"80001090" => n_pc <= X"80001094"; 
 n_reg10 <= X"00000000";

	when X"80001094" => 
 n_reg1 <= X"80001098"; n_pc <= reg18 + X"00000000";

	when X"80001098" => n_mem_addr <= reg2 + X"0000005c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"8000109C"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"8000109c" => n_mem_addr <= reg2 + X"00000058"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010A0"; n_reg8 <= (others => '0');n_reg8(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010a0" => n_mem_addr <= reg2 + X"00000054"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010A4"; n_reg9 <= (others => '0');n_reg9(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010a4" => n_mem_addr <= reg2 + X"00000050"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010A8"; n_reg18 <= (others => '0');n_reg18(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010a8" => n_mem_addr <= reg2 + X"0000004c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010AC"; n_reg19 <= (others => '0');n_reg19(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010ac" => n_mem_addr <= reg2 + X"00000048"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010B0"; n_reg20 <= (others => '0');n_reg20(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010b0" => n_mem_addr <= reg2 + X"00000044"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010B4"; n_reg21 <= (others => '0');n_reg21(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010b4" => n_mem_addr <= reg2 + X"00000040"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010B8"; n_reg22 <= (others => '0');n_reg22(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010b8" => n_mem_addr <= reg2 + X"0000003c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010BC"; n_reg23 <= (others => '0');n_reg23(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010bc" => n_mem_addr <= reg2 + X"00000038"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010C0"; n_reg24 <= (others => '0');n_reg24(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010c0" => n_mem_addr <= reg2 + X"00000034"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010C4"; n_reg25 <= (others => '0');n_reg25(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010c4" => n_mem_addr <= reg2 + X"00000030"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010C8"; n_reg26 <= (others => '0');n_reg26(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010c8" => n_pc <= X"800010cc"; 
 n_reg10 <= reg27;

	when X"800010cc" => n_mem_addr <= reg2 + X"0000002c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010D0"; n_reg27 <= (others => '0');n_reg27(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010d0" => n_pc <= X"800010d4"; 
 n_reg2 <= reg2 + X"00000060";

	when X"800010d4" => 
 n_pc <= reg1;

	when X"800010d8" => n_pc <= X"800010dc"; 
 n_reg15 <= reg23 + X"00000004";

	when X"800010dc" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000010"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then

 n_pc <= X"800010E0";
 end if;
	when X"800010e0" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010E4"; n_reg26 <= (others => '0');n_reg26(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800010e4" => n_pc <= X"800010e8"; 
 n_reg15 <= reg17;

	when X"800010e8" => n_pc <= X"800010ec"; 
 if signed(reg17) /= X"00000000" then n_pc <= X"800010f0"; end if;

	when X"800010ec" => n_pc <= X"800010f0"; 
 n_reg15 <= X"ffffffff";

	when X"800010f0" => n_pc <= X"800010f4"; 
 n_reg14 <= reg26 + reg15;

	when X"800010f4" => n_pc <= X"800010f8"; 
 n_reg15 <= reg26;

	when X"800010f8" => n_mem_addr <= reg15; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800010FC"; n_reg13 <= (others => '0');n_reg13(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"800010fc" => n_pc <= X"80001100"; 
 if signed(reg13) = X"00000000" then n_pc <= X"80001104"; end if;

	when X"80001100" => n_pc <= X"80001104"; 
 if signed(reg14) /= signed(reg15) then n_pc <= X"8000112c"; end if;

	when X"80001104" => n_pc <= X"80001108"; 
 n_reg23 <= reg6 and X"00000400";

	when X"80001108" => n_pc <= X"8000110c"; 
 n_reg25 <= reg15 - reg26;

	when X"8000110c" => n_pc <= X"80001110"; 
 if signed(reg23) = X"00000000" then n_pc <= X"80001118"; end if;

	when X"80001110" => n_pc <= X"80001114"; 
 if unsigned(reg17) >= unsigned(reg25) then n_pc <= X"80001118"; end if;

	when X"80001114" => n_pc <= X"80001118"; 
 n_reg25 <= reg17;

	when X"80001118" => n_pc <= X"8000111c"; 
 n_reg8 <= reg6 and X"00000002";

	when X"8000111c" => n_pc <= X"80001120"; 
 if signed(reg8) /= X"00000000" then n_pc <= X"80001184"; end if;

	when X"80001120" => n_pc <= X"80001124"; 
 n_reg12 <= reg27;

	when X"80001124" => n_pc <= X"80001128"; 
 n_reg6 <= reg25 - reg27;

	when X"80001128" => 
 n_pc <= X"80001164";

	when X"8000112c" => n_pc <= X"80001130"; 
 n_reg15 <= reg15 + X"00000001";

	when X"80001130" => 
 n_pc <= X"800010f8";

	when X"80001134" => n_pc <= X"80001138"; 
 n_reg14 <= reg12 + X"00000001";

	when X"80001138" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg6; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000113C";
 end if;
	when X"8000113c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000018"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001140";
 end if;
	when X"80001140" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000014"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001144";
 end if;
	when X"80001144" => n_pc <= X"80001148"; 
 n_reg13 <= reg19;

	when X"80001148" => n_pc <= X"8000114c"; 
 n_reg11 <= reg20;

	when X"8000114c" => n_pc <= X"80001150"; 
 n_reg10 <= X"00000020";

	when X"80001150" => 
 n_reg1 <= X"80001154"; n_pc <= reg18 + X"00000000";

	when X"80001154" => n_mem_addr <= reg2 + X"00000014"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001158"; n_reg14 <= (others => '0');n_reg14(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001158" => n_mem_addr <= reg2 + X"00000018"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"8000115C"; n_reg17 <= (others => '0');n_reg17(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"8000115c" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001160"; n_reg6 <= (others => '0');n_reg6(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001160" => n_pc <= X"80001164"; 
 n_reg12 <= reg14;

	when X"80001164" => n_pc <= X"80001168"; 
 n_reg14 <= reg12 + reg6;

	when X"80001168" => n_pc <= X"8000116c"; 
 if unsigned(reg14) < unsigned(reg24) then n_pc <= X"80001134"; end if;

	when X"8000116c" => n_pc <= X"80001170"; 
 n_reg14 <= X"00000000";

	when X"80001170" => n_pc <= X"80001174"; 
 if unsigned(reg24) < unsigned(reg25) then n_pc <= X"80001178"; end if;

	when X"80001174" => n_pc <= X"80001178"; 
 n_reg14 <= reg24 - reg25;

	when X"80001178" => n_pc <= X"8000117c"; 
 n_reg15 <= reg25 + X"00000001";

	when X"8000117c" => n_pc <= X"80001180"; 
 n_reg27 <= reg27 + reg14;

	when X"80001180" => n_pc <= X"80001184"; 
 n_reg25 <= reg14 + reg15;

	when X"80001184" => n_pc <= X"80001188"; 
 n_reg14 <= reg27;

	when X"80001188" => 
 n_pc <= X"800011b8";

	when X"8000118c" => n_pc <= X"80001190"; 
 n_reg17 <= reg13;

	when X"80001190" => n_pc <= X"80001194"; 
 n_reg6 <= reg14 + X"00000001";

	when X"80001194" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000018"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001198";
 end if;
	when X"80001198" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000014"; n_mem_wdata <= reg6; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000119C";
 end if;
	when X"8000119c" => n_pc <= X"800011a0"; 
 n_reg12 <= reg14;

	when X"800011a0" => n_pc <= X"800011a4"; 
 n_reg13 <= reg19;

	when X"800011a4" => n_pc <= X"800011a8"; 
 n_reg11 <= reg20;

	when X"800011a8" => 
 n_reg1 <= X"800011AC"; n_pc <= reg18 + X"00000000";

	when X"800011ac" => n_mem_addr <= reg2 + X"00000014"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800011B0"; n_reg6 <= (others => '0');n_reg6(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800011b0" => n_mem_addr <= reg2 + X"00000018"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800011B4"; n_reg17 <= (others => '0');n_reg17(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800011b4" => n_pc <= X"800011b8"; 
 n_reg14 <= reg6;

	when X"800011b8" => n_pc <= X"800011bc"; 
 n_reg13 <= reg14 - reg27;

	when X"800011bc" => n_pc <= X"800011c0"; 
 n_reg13 <= reg26 + reg13;

	when X"800011c0" => n_mem_addr <= reg13; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800011C4"; n_reg10 <= (others => '0');n_reg10(7 downto 0) <= mem_rdata(7 downto 0);
 end if;
	when X"800011c4" => n_pc <= X"800011c8"; 
 if signed(reg10) = X"00000000" then n_pc <= X"800011d4"; end if;

	when X"800011c8" => n_pc <= X"800011cc"; 
 if signed(reg23) = X"00000000" then n_pc <= X"80001190"; end if;

	when X"800011cc" => n_pc <= X"800011d0"; 
 n_reg13 <= reg17 + X"ffffffff";

	when X"800011d0" => n_pc <= X"800011d4"; 
 if signed(reg17) /= X"00000000" then n_pc <= X"8000118c"; end if;

	when X"800011d4" => n_pc <= X"800011d8"; 
 if signed(reg8) = X"00000000" then n_pc <= X"8000121c"; end if;

	when X"800011d8" => n_pc <= X"800011dc"; 
 n_reg12 <= reg14;

	when X"800011dc" => n_pc <= X"800011e0"; 
 n_reg8 <= reg25 - reg14;

	when X"800011e0" => 
 n_pc <= X"80001204";

	when X"800011e4" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000014"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800011E8";
 end if;
	when X"800011e8" => n_pc <= X"800011ec"; 
 n_reg13 <= reg19;

	when X"800011ec" => n_pc <= X"800011f0"; 
 n_reg11 <= reg20;

	when X"800011f0" => n_pc <= X"800011f4"; 
 n_reg10 <= X"00000020";

	when X"800011f4" => n_pc <= X"800011f8"; 
 n_reg23 <= reg12 + X"00000001";

	when X"800011f8" => 
 n_reg1 <= X"800011FC"; n_pc <= reg18 + X"00000000";

	when X"800011fc" => n_mem_addr <= reg2 + X"00000014"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001200"; n_reg14 <= (others => '0');n_reg14(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001200" => n_pc <= X"80001204"; 
 n_reg12 <= reg23;

	when X"80001204" => n_pc <= X"80001208"; 
 n_reg13 <= reg12 + reg8;

	when X"80001208" => n_pc <= X"8000120c"; 
 if unsigned(reg13) < unsigned(reg24) then n_pc <= X"800011e4"; end if;

	when X"8000120c" => n_pc <= X"80001210"; 
 n_reg13 <= X"00000000";

	when X"80001210" => n_pc <= X"80001214"; 
 if unsigned(reg24) < unsigned(reg25) then n_pc <= X"80001218"; end if;

	when X"80001214" => n_pc <= X"80001218"; 
 n_reg13 <= reg24 - reg25;

	when X"80001218" => n_pc <= X"8000121c"; 
 n_reg14 <= reg14 + reg13;

	when X"8000121c" => n_mem_addr <= reg2 + X"00000010"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001220"; n_reg23 <= (others => '0');n_reg23(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001220" => n_pc <= X"80001224"; 
 n_reg27 <= reg14;

	when X"80001224" => 
 n_pc <= X"80001074";

	when X"80001228" => n_pc <= X"8000122c"; 
 n_reg6 <= reg6 or X"00000021";

	when X"8000122c" => n_pc <= X"80001230"; 
 n_reg15 <= X"00000008";

	when X"80001230" => n_mem_addr <= reg23; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001234"; n_reg14 <= (others => '0');n_reg14(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001234" => n_pc <= X"80001238"; 
 n_reg8 <= reg23 + X"00000004";

	when X"80001238" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000004"; n_mem_wdata <= reg6; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000123C";
 end if;
	when X"8000123c" => mem_width <= "10"; n_mem_addr <= reg2; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001240";
 end if;
	when X"80001240" => n_pc <= X"80001244"; 
 n_reg16 <= X"00000010";

	when X"80001244" => 
 n_pc <= X"80000f90";

	when X"80001248" => n_pc <= X"8000124c"; 
 n_reg8 <= reg27 + X"00000001";

	when X"8000124c" => n_pc <= X"80001250"; 
 n_reg13 <= reg19;

	when X"80001250" => n_pc <= X"80001254"; 
 n_reg12 <= reg27;

	when X"80001254" => n_pc <= X"80001258"; 
 n_reg11 <= reg20;

	when X"80001258" => n_pc <= X"8000125c"; 
 n_reg10 <= X"00000025";

	when X"8000125c" => 
 n_reg1 <= X"80001260"; n_pc <= reg18 + X"00000000";

	when X"80001260" => n_pc <= X"80001264"; 
 n_reg27 <= reg8;

	when X"80001264" => 
 n_pc <= X"80001074";

	when X"80001268" => n_pc <= X"8000126c"; 
 n_reg16 <= X"00000008";

	when X"8000126c" => 
 n_pc <= X"80000ed4";

	when X"80001270" => n_pc <= X"80001274"; 
 n_reg16 <= X"00000002";

	when X"80001274" => 
 n_pc <= X"80000ed4";

	when X"80001278" => n_pc <= X"8000127c"; 
 n_reg2 <= reg2 + X"ffffffc0";

	when X"8000127c" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000002c"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001280";
 end if;
	when X"80001280" => n_pc <= X"80001284"; 
 n_reg13 <= reg10;

	when X"80001284" => n_pc <= X"80001288"; 
 n_reg10 <= X"80001000";

	when X"80001288" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000024"; n_mem_wdata <= reg11; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000128C";
 end if;
	when X"8000128c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000028"; n_mem_wdata <= reg12; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001290";
 end if;
	when X"80001290" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000030"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001294";
 end if;
	when X"80001294" => n_pc <= X"80001298"; 
 n_reg11 <= reg2 + X"00000008";

	when X"80001298" => n_pc <= X"8000129c"; 
 n_reg14 <= reg2 + X"00000024";

	when X"8000129c" => n_pc <= X"800012a0"; 
 n_reg12 <= X"ffffffff";

	when X"800012a0" => n_pc <= X"800012a4"; 
 n_reg10 <= reg10 + X"fffffbd4";

	when X"800012a4" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012A8";
 end if;
	when X"800012a8" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000034"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012AC";
 end if;
	when X"800012ac" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000038"; n_mem_wdata <= reg16; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012B0";
 end if;
	when X"800012b0" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012B4";
 end if;
	when X"800012b4" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012B8";
 end if;
	when X"800012b8" => 
 n_reg1 <= X"800012BC"; n_pc <= X"80000bf4";

	when X"800012bc" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800012C0"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800012c0" => n_pc <= X"800012c4"; 
 n_reg2 <= reg2 + X"00000040";

	when X"800012c4" => 
 n_pc <= reg1;

	when X"800012c8" => n_pc <= X"800012cc"; 
 n_reg2 <= reg2 + X"ffffffc0";

	when X"800012cc" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000002c"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012D0";
 end if;
	when X"800012d0" => n_pc <= X"800012d4"; 
 n_reg13 <= reg11;

	when X"800012d4" => n_pc <= X"800012d8"; 
 n_reg11 <= reg10;

	when X"800012d8" => n_pc <= X"800012dc"; 
 n_reg10 <= X"80001000";

	when X"800012dc" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000028"; n_mem_wdata <= reg12; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012E0";
 end if;
	when X"800012e0" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000030"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012E4";
 end if;
	when X"800012e4" => n_pc <= X"800012e8"; 
 n_reg12 <= X"ffffffff";

	when X"800012e8" => n_pc <= X"800012ec"; 
 n_reg14 <= reg2 + X"00000028";

	when X"800012ec" => n_pc <= X"800012f0"; 
 n_reg10 <= reg10 + X"fffff860";

	when X"800012f0" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012F4";
 end if;
	when X"800012f4" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000034"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012F8";
 end if;
	when X"800012f8" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000038"; n_mem_wdata <= reg16; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800012FC";
 end if;
	when X"800012fc" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001300";
 end if;
	when X"80001300" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001304";
 end if;
	when X"80001304" => 
 n_reg1 <= X"80001308"; n_pc <= X"80000bf4";

	when X"80001308" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"8000130C"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"8000130c" => n_pc <= X"80001310"; 
 n_reg2 <= reg2 + X"00000040";

	when X"80001310" => 
 n_pc <= reg1;

	when X"80001314" => n_pc <= X"80001318"; 
 n_reg2 <= reg2 + X"ffffffc0";

	when X"80001318" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000002c"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000131C";
 end if;
	when X"8000131c" => n_pc <= X"80001320"; 
 n_reg13 <= reg12;

	when X"80001320" => n_pc <= X"80001324"; 
 n_reg12 <= reg11;

	when X"80001324" => n_pc <= X"80001328"; 
 n_reg11 <= reg10;

	when X"80001328" => n_pc <= X"8000132c"; 
 n_reg10 <= X"80001000";

	when X"8000132c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000030"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001330";
 end if;
	when X"80001330" => n_pc <= X"80001334"; 
 n_reg10 <= reg10 + X"fffff860";

	when X"80001334" => n_pc <= X"80001338"; 
 n_reg14 <= reg2 + X"0000002c";

	when X"80001338" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000133C";
 end if;
	when X"8000133c" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000034"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001340";
 end if;
	when X"80001340" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000038"; n_mem_wdata <= reg16; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001344";
 end if;
	when X"80001344" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"80001348";
 end if;
	when X"80001348" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000134C";
 end if;
	when X"8000134c" => 
 n_reg1 <= X"80001350"; n_pc <= X"80000bf4";

	when X"80001350" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001354"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001354" => n_pc <= X"80001358"; 
 n_reg2 <= reg2 + X"00000040";

	when X"80001358" => 
 n_pc <= reg1;

	when X"8000135c" => n_pc <= X"80001360"; 
 n_reg2 <= reg2 + X"ffffffe0";

	when X"80001360" => n_pc <= X"80001364"; 
 n_reg13 <= reg10;

	when X"80001364" => n_pc <= X"80001368"; 
 n_reg10 <= X"80001000";

	when X"80001368" => n_pc <= X"8000136c"; 
 n_reg14 <= reg11;

	when X"8000136c" => n_pc <= X"80001370"; 
 n_reg12 <= X"ffffffff";

	when X"80001370" => n_pc <= X"80001374"; 
 n_reg11 <= reg2 + X"0000000c";

	when X"80001374" => n_pc <= X"80001378"; 
 n_reg10 <= reg10 + X"fffffbd4";

	when X"80001378" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"8000137C";
 end if;
	when X"8000137c" => 
 n_reg1 <= X"80001380"; n_pc <= X"80000bf4";

	when X"80001380" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"80001384"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"80001384" => n_pc <= X"80001388"; 
 n_reg2 <= reg2 + X"00000020";

	when X"80001388" => 
 n_pc <= reg1;

	when X"8000138c" => n_pc <= X"80001390"; 
 n_reg14 <= reg13;

	when X"80001390" => n_pc <= X"80001394"; 
 n_reg13 <= reg12;

	when X"80001394" => n_pc <= X"80001398"; 
 n_reg12 <= reg11;

	when X"80001398" => n_pc <= X"8000139c"; 
 n_reg11 <= reg10;

	when X"8000139c" => n_pc <= X"800013a0"; 
 n_reg10 <= X"80001000";

	when X"800013a0" => n_pc <= X"800013a4"; 
 n_reg10 <= reg10 + X"fffff860";

	when X"800013a4" => 
 n_pc <= X"80000bf4";

	when X"800013a8" => n_pc <= X"800013ac"; 
 n_reg2 <= reg2 + X"ffffffc0";

	when X"800013ac" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000008"; n_mem_wdata <= reg10; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013B0";
 end if;
	when X"800013b0" => n_pc <= X"800013b4"; 
 n_reg10 <= X"80001000";

	when X"800013b4" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000002c"; n_mem_wdata <= reg13; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013B8";
 end if;
	when X"800013b8" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000030"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013BC";
 end if;
	when X"800013bc" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000000c"; n_mem_wdata <= reg11; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013C0";
 end if;
	when X"800013c0" => n_pc <= X"800013c4"; 
 n_reg14 <= reg2 + X"0000002c";

	when X"800013c4" => n_pc <= X"800013c8"; 
 n_reg13 <= reg12;

	when X"800013c8" => n_pc <= X"800013cc"; 
 n_reg11 <= reg2 + X"00000008";

	when X"800013cc" => n_pc <= X"800013d0"; 
 n_reg12 <= X"ffffffff";

	when X"800013d0" => n_pc <= X"800013d4"; 
 n_reg10 <= reg10 + X"fffffbe0";

	when X"800013d4" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000001c"; n_mem_wdata <= reg1; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013D8";
 end if;
	when X"800013d8" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000034"; n_mem_wdata <= reg15; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013DC";
 end if;
	when X"800013dc" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000038"; n_mem_wdata <= reg16; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013E0";
 end if;
	when X"800013e0" => mem_width <= "10"; n_mem_addr <= reg2 + X"0000003c"; n_mem_wdata <= reg17; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013E4";
 end if;
	when X"800013e4" => mem_width <= "10"; n_mem_addr <= reg2 + X"00000004"; n_mem_wdata <= reg14; mem_we <= '1'; if mem_wack = '1' then
 n_pc <= X"800013E8";
 end if;
	when X"800013e8" => 
 n_reg1 <= X"800013EC"; n_pc <= X"80000bf4";

	when X"800013ec" => n_mem_addr <= reg2 + X"0000001c"; mem_re <= '1'; if mem_rdy = '1' then
 n_pc <= X"800013F0"; n_reg1 <= (others => '0');n_reg1(31 downto 0) <= mem_rdata(31 downto 0);
 end if;
	when X"800013f0" => n_pc <= X"800013f4"; 
 n_reg2 <= reg2 + X"00000040";

	when X"800013f4" => 
 n_pc <= reg1;

	when X"800013f8" =>
		
	when others =>
		n_pc <= X"800013f8";
end case;
end process;

end Behavioural;